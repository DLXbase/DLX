package alu_type is
	type aluOp is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, FUNCRSL, FUNCRR, SGE, SLE, SNE, aluNOP);
end alu_type;
