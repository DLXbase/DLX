package alu_type is
	type aluOp is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, FUNCRL, FUNCRR, SGE, SLE, SNE, NOP);
end alu_type;
